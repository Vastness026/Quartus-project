library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LEDcount_down is
port (
		clk : in std_logic;
		reset : in std_logic;
		rows : out std_logic_vector(7 downto 0);
		cols  : out std_logic_vector(7 downto 0);
		lose : out std_logic := '0'
);
end LEDcount_down;

architecture oo of LEDcount_down is
	
	signal clk_counter : integer := 0;
	signal matrix_counter : integer := 30;
	signal row_counter : unsigned(2 downto 0);

	type matrix_type is array (0 to 7) of std_logic_vector(7 downto 0);
	type matrix_array is array(0 to 30) of matrix_type;
	
	signal matrix3d : matrix_array;
	
	
	
begin

	matrix3d(0) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','0','0','1','1','0'),
	('1','0','0','1','1','0','0','1'),
	('1','0','0','1','1','0','0','1'),
	('1','0','0','1','1','0','0','1'),
	('0','1','1','0','0','1','1','0'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(1) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','0','0','0','1','0'),
	('1','0','0','1','0','0','1','0'),
	('1','0','0','1','0','0','1','0'),
	('1','0','0','1','0','0','1','0'),
	('0','1','1','0','0','0','1','0'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(2) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','0','0','1','1','1'),
	('1','0','0','1','0','0','0','1'),
	('1','0','0','1','0','1','1','1'),
	('1','0','0','1','0','1','0','0'),
	('0','1','1','0','0','1','1','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(3) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','0','0','1','1','1'),
	('1','0','0','1','0','0','0','1'),
	('1','0','0','1','0','1','1','1'),
	('1','0','0','1','0','0','0','1'),
	('0','1','1','0','0','1','1','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(4) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','0','0','1','0','1'),
	('1','0','0','1','0','1','0','1'),
	('1','0','0','1','0','1','1','1'),
	('1','0','0','1','0','0','0','1'),
	('0','1','1','0','0','0','0','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(5) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','0','0','1','1','1'),
	('1','0','0','1','0','1','0','0'),
	('1','0','0','1','0','1','1','1'),
	('1','0','0','1','0','0','0','1'),
	('0','1','1','0','0','1','1','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(6) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','0','0','1','1','1'),
	('1','0','0','1','0','1','0','0'),
	('1','0','0','1','0','1','1','1'),
	('1','0','0','1','0','1','0','1'),
	('0','1','1','0','0','1','1','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(7) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','0','0','1','1','1'),
	('1','0','0','1','0','1','0','1'),
	('1','0','0','1','0','1','0','1'),
	('1','0','0','1','0','0','0','1'),
	('0','1','1','0','0','0','0','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(8) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','0','0','1','1','1'),
	('1','0','0','1','0','1','0','1'),
	('1','0','0','1','0','1','1','1'),
	('1','0','0','1','0','1','0','1'),
	('0','1','1','0','0','1','1','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(9) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','0','0','1','1','1'),
	('1','0','0','1','0','1','0','1'),
	('1','0','0','1','0','1','1','1'),
	('1','0','0','1','0','0','0','1'),
	('0','1','1','0','0','0','0','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(10) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','0','1','0','0','1','1','0'),
	('0','0','1','0','1','0','0','1'),
	('0','0','1','0','1','0','0','1'),
	('0','0','1','0','1','0','0','1'),
	('0','0','1','0','0','1','1','0'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(11) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','0','1','0','0','0','1','0'),
	('0','0','1','0','0','0','1','0'),
	('0','0','1','0','0','0','1','0'),
	('0','0','1','0','0','0','1','0'),
	('0','0','1','0','0','0','1','0'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(12) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','0','1','0','0','1','1','1'),
	('0','0','1','0','0','0','0','1'),
	('0','0','1','0','0','1','1','1'),
	('0','0','1','0','0','1','0','0'),
	('0','0','1','0','0','1','1','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(13) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','0','1','0','0','1','1','1'),
	('0','0','1','0','0','0','0','1'),
	('0','0','1','0','0','1','1','1'),
	('0','0','1','0','0','0','0','1'),
	('0','0','1','0','0','1','1','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(14) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','0','1','0','0','1','0','1'),
	('0','0','1','0','0','1','0','1'),
	('0','0','1','0','0','1','1','1'),
	('0','0','1','0','0','0','0','1'),
	('0','0','1','0','0','0','0','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(15) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','0','1','0','0','1','1','1'),
	('0','0','1','0','0','1','0','0'),
	('0','0','1','0','0','1','1','1'),
	('0','0','1','0','0','0','0','1'),
	('0','0','1','0','0','1','1','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(16) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','0','1','0','0','1','1','1'),
	('0','0','1','0','0','1','0','0'),
	('0','0','1','0','0','1','1','1'),
	('0','0','1','0','0','1','0','1'),
	('0','0','1','0','0','1','1','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(17) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','0','1','0','0','1','1','1'),
	('0','0','1','0','0','1','0','1'),
	('0','0','1','0','0','1','0','1'),
	('0','0','1','0','0','0','0','1'),
	('0','0','1','0','0','0','0','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(18) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','0','1','0','0','1','1','1'),
	('0','0','1','0','0','1','0','1'),
	('0','0','1','0','0','1','1','1'),
	('0','0','1','0','0','1','0','1'),
	('0','0','1','0','0','1','1','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(19) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','0','1','0','0','1','1','1'),
	('0','0','1','0','0','1','0','1'),
	('0','0','1','0','0','1','1','1'),
	('0','0','1','0','0','0','0','1'),
	('0','0','1','0','0','0','0','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(20) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','1','0','1','1','0'),
	('0','0','0','1','1','0','0','1'),
	('0','1','1','1','1','0','0','1'),
	('0','1','0','0','1','0','0','1'),
	('0','1','1','1','0','1','1','0'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(21) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','1','0','0','1','0'),
	('0','0','0','1','0','0','1','0'),
	('0','1','1','1','0','0','1','0'),
	('0','1','0','0','0','0','1','0'),
	('0','1','1','1','0','0','1','0'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(22) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','1','0','1','1','1'),
	('0','0','0','1','0','0','0','1'),
	('0','1','1','1','0','1','1','1'),
	('0','1','0','0','0','1','0','0'),
	('0','1','1','1','0','1','1','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(23) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','1','0','1','1','1'),
	('0','0','0','1','0','0','0','1'),
	('0','1','1','1','0','1','1','1'),
	('0','1','0','0','0','0','0','1'),
	('0','1','1','1','0','1','1','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(24) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','1','0','1','0','1'),
	('0','0','0','1','0','1','0','1'),
	('0','1','1','1','0','1','1','1'),
	('0','1','0','0','0','0','0','1'),
	('0','1','1','1','0','0','0','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(25) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','1','0','1','1','1'),
	('0','0','0','1','0','1','0','0'),
	('0','1','1','1','0','1','1','1'),
	('0','1','0','0','0','0','0','1'),
	('0','1','1','1','0','1','1','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(26) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','1','0','1','1','1'),
	('0','0','0','1','0','1','0','0'),
	('0','1','1','1','0','1','1','1'),
	('0','1','0','0','0','1','0','1'),
	('0','1','1','1','0','1','1','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(27) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','1','0','1','1','1'),
	('0','0','0','1','0','1','0','1'),
	('0','1','1','1','0','1','0','1'),
	('0','1','0','0','0','0','0','1'),
	('0','1','1','1','0','0','0','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(28) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','1','0','1','1','1'),
	('0','0','0','1','0','1','0','1'),
	('0','1','1','1','0','1','1','1'),
	('0','1','0','0','0','1','0','1'),
	('0','1','1','1','0','1','1','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(29) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','1','0','1','1','1'),
	('0','0','0','1','0','1','0','1'),
	('0','1','1','1','0','1','1','1'),
	('0','1','0','0','0','0','0','1'),
	('0','1','1','1','0','0','0','1'),
	('0','0','0','0','0','0','0','0')
	);
	matrix3d(30) <= (
	('0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0'),
	('0','1','1','1','0','1','1','0'),
	('0','0','0','1','1','0','0','1'),
	('0','1','1','1','1','0','0','1'),
	('0','0','0','1','1','0','0','1'),
	('0','1','1','1','0','1','1','0'),
	('0','0','0','0','0','0','0','0')
	);
	COUNTER_PROC : process(clk)
	begin
		if reset = '0' then
		
			if rising_edge(clk) then
		
				if (clk_counter > 10 or clk_counter = 10) then
			
					clk_counter <= 0;
					if matrix_counter > 0 then
						matrix_counter <= matrix_counter - 1;
					end if;
				
				else
					clk_counter <= clk_counter + 1;
				end if;
				
				if matrix_counter > 0 then
					row_counter <= row_counter + 1;
				end if;
				
			end if;
			
		else
			clk_counter <= 0;
			matrix_counter <= 30;
		end if;
	end process;
	
	OUTPUT_PROC : process(row_counter)
	begin
		
		cols <= matrix3d(matrix_counter)(to_integer(row_counter));
		
		rows <= (others => '0');
		rows(to_integer(row_counter)) <= '1';
		
		if reset = '1' then
			rows <= (others => '0');
			cols <= (others => '0');
		end if;
		
		if matrix_counter = 0 then
			lose <= '1';
			rows <= (others => '0');
			cols <= (others => '0');
		else
			lose <= '0';
		end if;
		
	end process;
	
end architecture;
	